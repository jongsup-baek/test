mdoule
\endmodule
